library IEEE;
use IEEE.std_logic_1164.all;

package testbench_pkg is
   constant FILE_NAME : string := "chk_sim_sig_advanced.txt";

   constant N_TEST_WORDS : integer := 1642; 
   type t_test_words     is array (1 to N_TEST_WORDS) 
                                  of string(1 to 15);
   constant test_words : t_test_words :=
   ( 
     "067108088#     ",
     "167108088#     ",
     "267108088#     ",
     "367108088#     ",
     "467108088#     ",
     "567108088#     ",
     "667108088#     ",
     "767108088#     ",
     "867108088#     ",
     "967108088#     ",
     "A67108088#     ",
     "B67108088#     ",
     "C67108088#     ",
     "D67108088#     ",
     "*67108088#     ",
     "707108088#     ",
     "717108088#     ",
     "727108088#     ",
     "737108088#     ",
     "747108088#     ",
     "757108088#     ",
     "767108088#     ",
     "777108088#     ",
     "787108088#     ",
     "797108088#     ",
     "7A7108088#     ",
     "7B7108088#     ",
     "7C7108088#     ",
     "7D7108088#     ",
     "7*7108088#     ",
     "760108088#     ",
     "761108088#     ",
     "762108088#     ",
     "763108088#     ",
     "764108088#     ",
     "765108088#     ",
     "766108088#     ",
     "767108088#     ",
     "768108088#     ",
     "769108088#     ",
     "76A108088#     ",
     "76B108088#     ",
     "76C108088#     ",
     "76D108088#     ",
     "76*108088#     ",
     "767008088#     ",
     "767108088#     ",
     "767208088#     ",
     "767308088#     ",
     "767408088#     ",
     "767508088#     ",
     "767608088#     ",
     "767708088#     ",
     "767808088#     ",
     "767908088#     ",
     "767A08088#     ",
     "767B08088#     ",
     "767C08088#     ",
     "767D08088#     ",
     "767*08088#     ",
     "767108088#     ",
     "767118088#     ",
     "767128088#     ",
     "767138088#     ",
     "767148088#     ",
     "767158088#     ",
     "767168088#     ",
     "767178088#     ",
     "767188088#     ",
     "767198088#     ",
     "7671A8088#     ",
     "7671B8088#     ",
     "7671C8088#     ",
     "7671D8088#     ",
     "7671*8088#     ",
     "767100088#     ",
     "767101088#     ",
     "767102088#     ",
     "767103088#     ",
     "767104088#     ",
     "767105088#     ",
     "767106088#     ",
     "767107088#     ",
     "767108088#     ",
     "767109088#     ",
     "76710A088#     ",
     "76710B088#     ",
     "76710C088#     ",
     "76710D088#     ",
     "76710*088#     ",
     "767108088#     ",
     "767108188#     ",
     "767108288#     ",
     "767108388#     ",
     "767108488#     ",
     "767108588#     ",
     "767108688#     ",
     "767108788#     ",
     "767108888#     ",
     "767108988#     ",
     "767108A88#     ",
     "767108B88#     ",
     "767108C88#     ",
     "767108D88#     ",
     "767108*88#     ",
     "767108008#     ",
     "767108018#     ",
     "767108028#     ",
     "767108038#     ",
     "767108048#     ",
     "767108058#     ",
     "767108068#     ",
     "767108078#     ",
     "767108088#     ",
     "767108098#     ",
     "7671080A8#     ",
     "7671080B8#     ",
     "7671080C8#     ",
     "7671080D8#     ",
     "7671080*8#     ",
     "767108080#     ",
     "767108081#     ",
     "767108082#     ",
     "767108083#     ",
     "767108084#     ",
     "767108085#     ",
     "767108086#     ",
     "767108087#     ",
     "767108088#     ",
     "767108089#     ",
     "76710808A#     ",
     "76710808B#     ",
     "76710808C#     ",
     "76710808D#     ",
     "76710808*#     ",
     "00#            ",
     "01#            ",
     "02#            ",
     "03#            ",
     "04#            ",
     "05#            ",
     "06#            ",
     "07#            ",
     "08#            ",
     "09#            ",
     "0A#            ",
     "0B#            ",
     "0C#            ",
     "0D#            ",
     "0*#            ",
     "0#             ",
     "10#            ",
     "11#            ",
     "12#            ",
     "13#            ",
     "14#            ",
     "15#            ",
     "16#            ",
     "17#            ",
     "18#            ",
     "19#            ",
     "1A#            ",
     "1B#            ",
     "1C#            ",
     "1D#            ",
     "1*#            ",
     "1#             ",
     "20#            ",
     "21#            ",
     "22#            ",
     "23#            ",
     "24#            ",
     "25#            ",
     "26#            ",
     "27#            ",
     "28#            ",
     "29#            ",
     "2A#            ",
     "2B#            ",
     "2C#            ",
     "2D#            ",
     "2*#            ",
     "2#             ",
     "30#            ",
     "31#            ",
     "32#            ",
     "33#            ",
     "34#            ",
     "35#            ",
     "36#            ",
     "37#            ",
     "38#            ",
     "39#            ",
     "3A#            ",
     "3B#            ",
     "3C#            ",
     "3D#            ",
     "3*#            ",
     "3#             ",
     "40#            ",
     "41#            ",
     "42#            ",
     "43#            ",
     "44#            ",
     "45#            ",
     "46#            ",
     "47#            ",
     "48#            ",
     "49#            ",
     "4A#            ",
     "4B#            ",
     "4C#            ",
     "4D#            ",
     "4*#            ",
     "4#             ",
     "50#            ",
     "51#            ",
     "52#            ",
     "53#            ",
     "54#            ",
     "55#            ",
     "56#            ",
     "57#            ",
     "58#            ",
     "59#            ",
     "5A#            ",
     "5B#            ",
     "5C#            ",
     "5D#            ",
     "5*#            ",
     "5#             ",
     "60#            ",
     "61#            ",
     "62#            ",
     "63#            ",
     "64#            ",
     "65#            ",
     "66#            ",
     "67#            ",
     "68#            ",
     "69#            ",
     "6A#            ",
     "6B#            ",
     "6C#            ",
     "6D#            ",
     "6*#            ",
     "6#             ",
     "70#            ",
     "71#            ",
     "72#            ",
     "73#            ",
     "74#            ",
     "75#            ",
     "76#            ",
     "77#            ",
     "78#            ",
     "79#            ",
     "7A#            ",
     "7B#            ",
     "7C#            ",
     "7D#            ",
     "7*#            ",
     "7#             ",
     "80#            ",
     "81#            ",
     "82#            ",
     "83#            ",
     "84#            ",
     "85#            ",
     "86#            ",
     "87#            ",
     "88#            ",
     "89#            ",
     "8A#            ",
     "8B#            ",
     "8C#            ",
     "8D#            ",
     "8*#            ",
     "8#             ",
     "90#            ",
     "91#            ",
     "92#            ",
     "93#            ",
     "94#            ",
     "95#            ",
     "96#            ",
     "97#            ",
     "98#            ",
     "99#            ",
     "9A#            ",
     "9B#            ",
     "9C#            ",
     "9D#            ",
     "9*#            ",
     "9#             ",
     "A0#            ",
     "A1#            ",
     "A2#            ",
     "A3#            ",
     "A4#            ",
     "A5#            ",
     "A6#            ",
     "A7#            ",
     "A8#            ",
     "A9#            ",
     "AA#            ",
     "AB#            ",
     "AC#            ",
     "AD#            ",
     "A*#            ",
     "A#             ",
     "B0#            ",
     "B1#            ",
     "B2#            ",
     "B3#            ",
     "B4#            ",
     "B5#            ",
     "B6#            ",
     "B7#            ",
     "B8#            ",
     "B9#            ",
     "BA#            ",
     "BB#            ",
     "BC#            ",
     "BD#            ",
     "B*#            ",
     "B#             ",
     "C0#            ",
     "C1#            ",
     "C2#            ",
     "C3#            ",
     "C4#            ",
     "C5#            ",
     "C6#            ",
     "C7#            ",
     "C8#            ",
     "C9#            ",
     "CA#            ",
     "CB#            ",
     "CC#            ",
     "CD#            ",
     "C*#            ",
     "C#             ",
     "D0#            ",
     "D1#            ",
     "D2#            ",
     "D3#            ",
     "D4#            ",
     "D5#            ",
     "D6#            ",
     "D7#            ",
     "D8#            ",
     "D9#            ",
     "DA#            ",
     "DB#            ",
     "DC#            ",
     "DD#            ",
     "D*#            ",
     "D#             ",
     "*0#            ",
     "*1#            ",
     "*2#            ",
     "*3#            ",
     "*4#            ",
     "*5#            ",
     "*6#            ",
     "*7#            ",
     "*8#            ",
     "*9#            ",
     "*A#            ",
     "*B#            ",
     "*C#            ",
     "*D#            ",
     "**#            ",
     "*#             ",
     "767108000#     ",
     "767108001#     ",
     "767108002#     ",
     "767108003#     ",
     "767108004#     ",
     "767108005#     ",
     "767108006#     ",
     "767108007#     ",
     "767108008#     ",
     "767108009#     ",
     "76710800A#     ",
     "76710800B#     ",
     "76710800C#     ",
     "76710800D#     ",
     "76710800*#     ",
     "76710800#      ",
     "767108010#     ",
     "767108011#     ",
     "767108012#     ",
     "767108013#     ",
     "767108014#     ",
     "767108015#     ",
     "767108016#     ",
     "767108017#     ",
     "767108018#     ",
     "767108019#     ",
     "76710801A#     ",
     "76710801B#     ",
     "76710801C#     ",
     "76710801D#     ",
     "76710801*#     ",
     "76710801#      ",
     "767108020#     ",
     "767108021#     ",
     "767108022#     ",
     "767108023#     ",
     "767108024#     ",
     "767108025#     ",
     "767108026#     ",
     "767108027#     ",
     "767108028#     ",
     "767108029#     ",
     "76710802A#     ",
     "76710802B#     ",
     "76710802C#     ",
     "76710802D#     ",
     "76710802*#     ",
     "76710802#      ",
     "767108030#     ",
     "767108031#     ",
     "767108032#     ",
     "767108033#     ",
     "767108034#     ",
     "767108035#     ",
     "767108036#     ",
     "767108037#     ",
     "767108038#     ",
     "767108039#     ",
     "76710803A#     ",
     "76710803B#     ",
     "76710803C#     ",
     "76710803D#     ",
     "76710803*#     ",
     "76710803#      ",
     "767108040#     ",
     "767108041#     ",
     "767108042#     ",
     "767108043#     ",
     "767108044#     ",
     "767108045#     ",
     "767108046#     ",
     "767108047#     ",
     "767108048#     ",
     "767108049#     ",
     "76710804A#     ",
     "76710804B#     ",
     "76710804C#     ",
     "76710804D#     ",
     "76710804*#     ",
     "76710804#      ",
     "767108050#     ",
     "767108051#     ",
     "767108052#     ",
     "767108053#     ",
     "767108054#     ",
     "767108055#     ",
     "767108056#     ",
     "767108057#     ",
     "767108058#     ",
     "767108059#     ",
     "76710805A#     ",
     "76710805B#     ",
     "76710805C#     ",
     "76710805D#     ",
     "76710805*#     ",
     "76710805#      ",
     "767108060#     ",
     "767108061#     ",
     "767108062#     ",
     "767108063#     ",
     "767108064#     ",
     "767108065#     ",
     "767108066#     ",
     "767108067#     ",
     "767108068#     ",
     "767108069#     ",
     "76710806A#     ",
     "76710806B#     ",
     "76710806C#     ",
     "76710806D#     ",
     "76710806*#     ",
     "76710806#      ",
     "767108070#     ",
     "767108071#     ",
     "767108072#     ",
     "767108073#     ",
     "767108074#     ",
     "767108075#     ",
     "767108076#     ",
     "767108077#     ",
     "767108078#     ",
     "767108079#     ",
     "76710807A#     ",
     "76710807B#     ",
     "76710807C#     ",
     "76710807D#     ",
     "76710807*#     ",
     "76710807#      ",
     "767108080#     ",
     "767108081#     ",
     "767108082#     ",
     "767108083#     ",
     "767108084#     ",
     "767108085#     ",
     "767108086#     ",
     "767108087#     ",
     "767108088#     ",
     "767108089#     ",
     "76710808A#     ",
     "76710808B#     ",
     "76710808C#     ",
     "76710808D#     ",
     "76710808*#     ",
     "76710808#      ",
     "767108090#     ",
     "767108091#     ",
     "767108092#     ",
     "767108093#     ",
     "767108094#     ",
     "767108095#     ",
     "767108096#     ",
     "767108097#     ",
     "767108098#     ",
     "767108099#     ",
     "76710809A#     ",
     "76710809B#     ",
     "76710809C#     ",
     "76710809D#     ",
     "76710809*#     ",
     "76710809#      ",
     "7671080A0#     ",
     "7671080A1#     ",
     "7671080A2#     ",
     "7671080A3#     ",
     "7671080A4#     ",
     "7671080A5#     ",
     "7671080A6#     ",
     "7671080A7#     ",
     "7671080A8#     ",
     "7671080A9#     ",
     "7671080AA#     ",
     "7671080AB#     ",
     "7671080AC#     ",
     "7671080AD#     ",
     "7671080A*#     ",
     "7671080A#      ",
     "7671080B0#     ",
     "7671080B1#     ",
     "7671080B2#     ",
     "7671080B3#     ",
     "7671080B4#     ",
     "7671080B5#     ",
     "7671080B6#     ",
     "7671080B7#     ",
     "7671080B8#     ",
     "7671080B9#     ",
     "7671080BA#     ",
     "7671080BB#     ",
     "7671080BC#     ",
     "7671080BD#     ",
     "7671080B*#     ",
     "7671080B#      ",
     "7671080C0#     ",
     "7671080C1#     ",
     "7671080C2#     ",
     "7671080C3#     ",
     "7671080C4#     ",
     "7671080C5#     ",
     "7671080C6#     ",
     "7671080C7#     ",
     "7671080C8#     ",
     "7671080C9#     ",
     "7671080CA#     ",
     "7671080CB#     ",
     "7671080CC#     ",
     "7671080CD#     ",
     "7671080C*#     ",
     "7671080C#      ",
     "7671080D0#     ",
     "7671080D1#     ",
     "7671080D2#     ",
     "7671080D3#     ",
     "7671080D4#     ",
     "7671080D5#     ",
     "7671080D6#     ",
     "7671080D7#     ",
     "7671080D8#     ",
     "7671080D9#     ",
     "7671080DA#     ",
     "7671080DB#     ",
     "7671080DC#     ",
     "7671080DD#     ",
     "7671080D*#     ",
     "7671080D#      ",
     "7671080*0#     ",
     "7671080*1#     ",
     "7671080*2#     ",
     "7671080*3#     ",
     "7671080*4#     ",
     "7671080*5#     ",
     "7671080*6#     ",
     "7671080*7#     ",
     "7671080*8#     ",
     "7671080*9#     ",
     "7671080*A#     ",
     "7671080*B#     ",
     "7671080*C#     ",
     "7671080*D#     ",
     "7671080**#     ",
     "7671080*#      ",
     "0767108088#    ",
     "1767108088#    ",
     "2767108088#    ",
     "3767108088#    ",
     "4767108088#    ",
     "5767108088#    ",
     "6767108088#    ",
     "7767108088#    ",
     "8767108088#    ",
     "9767108088#    ",
     "A767108088#    ",
     "B767108088#    ",
     "C767108088#    ",
     "D767108088#    ",
     "*767108088#    ",
     "7067108088#    ",
     "7167108088#    ",
     "7267108088#    ",
     "7367108088#    ",
     "7467108088#    ",
     "7567108088#    ",
     "7667108088#    ",
     "7767108088#    ",
     "7867108088#    ",
     "7967108088#    ",
     "7A67108088#    ",
     "7B67108088#    ",
     "7C67108088#    ",
     "7D67108088#    ",
     "7*67108088#    ",
     "7607108088#    ",
     "7617108088#    ",
     "7627108088#    ",
     "7637108088#    ",
     "7647108088#    ",
     "7657108088#    ",
     "7667108088#    ",
     "7677108088#    ",
     "7687108088#    ",
     "7697108088#    ",
     "76A7108088#    ",
     "76B7108088#    ",
     "76C7108088#    ",
     "76D7108088#    ",
     "76*7108088#    ",
     "7670108088#    ",
     "7671108088#    ",
     "7672108088#    ",
     "7673108088#    ",
     "7674108088#    ",
     "7675108088#    ",
     "7676108088#    ",
     "7677108088#    ",
     "7678108088#    ",
     "7679108088#    ",
     "767A108088#    ",
     "767B108088#    ",
     "767C108088#    ",
     "767D108088#    ",
     "767*108088#    ",
     "7671008088#    ",
     "7671108088#    ",
     "7671208088#    ",
     "7671308088#    ",
     "7671408088#    ",
     "7671508088#    ",
     "7671608088#    ",
     "7671708088#    ",
     "7671808088#    ",
     "7671908088#    ",
     "7671A08088#    ",
     "7671B08088#    ",
     "7671C08088#    ",
     "7671D08088#    ",
     "7671*08088#    ",
     "7671008088#    ",
     "7671018088#    ",
     "7671028088#    ",
     "7671038088#    ",
     "7671048088#    ",
     "7671058088#    ",
     "7671068088#    ",
     "7671078088#    ",
     "7671088088#    ",
     "7671098088#    ",
     "76710A8088#    ",
     "76710B8088#    ",
     "76710C8088#    ",
     "76710D8088#    ",
     "76710*8088#    ",
     "7671080088#    ",
     "7671081088#    ",
     "7671082088#    ",
     "7671083088#    ",
     "7671084088#    ",
     "7671085088#    ",
     "7671086088#    ",
     "7671087088#    ",
     "7671088088#    ",
     "7671089088#    ",
     "767108A088#    ",
     "767108B088#    ",
     "767108C088#    ",
     "767108D088#    ",
     "767108*088#    ",
     "7671080088#    ",
     "7671080188#    ",
     "7671080288#    ",
     "7671080388#    ",
     "7671080488#    ",
     "7671080588#    ",
     "7671080688#    ",
     "7671080788#    ",
     "7671080888#    ",
     "7671080988#    ",
     "7671080A88#    ",
     "7671080B88#    ",
     "7671080C88#    ",
     "7671080D88#    ",
     "7671080*88#    ",
     "7671080808#    ",
     "7671080818#    ",
     "7671080828#    ",
     "7671080838#    ",
     "7671080848#    ",
     "7671080858#    ",
     "7671080868#    ",
     "7671080878#    ",
     "7671080888#    ",
     "7671080898#    ",
     "76710808A8#    ",
     "76710808B8#    ",
     "76710808C8#    ",
     "76710808D8#    ",
     "76710808*8#    ",
     "7671080880#    ",
     "7671080881#    ",
     "7671080882#    ",
     "7671080883#    ",
     "7671080884#    ",
     "7671080885#    ",
     "7671080886#    ",
     "7671080887#    ",
     "7671080888#    ",
     "7671080889#    ",
     "767108088A#    ",
     "767108088B#    ",
     "767108088C#    ",
     "767108088D#    ",
     "767108088*#    ",
     "67108088#      ",
     "77108088#      ",
     "76108088#      ",
     "76708088#      ",
     "76718088#      ",
     "76710088#      ",
     "76710888#      ",
     "76710808#      ",
     "76710808#      ",
     "#              ",
     "7#             ",
     "76#            ",
     "767#           ",
     "7671#          ",
     "76710#         ",
     "767108#        ",
     "7671080#       ",
     "76710808#      ",
     "767108088#     ",
     "767108088#     ",
     "67108088#      ",
     "7108088#       ",
     "108088#        ",
     "08088#         ",
     "8088#          ",
     "088#           ",
     "88#            ",
     "8#             ",
     "#              ",
     "0671216177#    ",
     "1671216177#    ",
     "2671216177#    ",
     "3671216177#    ",
     "4671216177#    ",
     "5671216177#    ",
     "6671216177#    ",
     "7671216177#    ",
     "8671216177#    ",
     "9671216177#    ",
     "A671216177#    ",
     "B671216177#    ",
     "C671216177#    ",
     "D671216177#    ",
     "*671216177#    ",
     "7071216177#    ",
     "7171216177#    ",
     "7271216177#    ",
     "7371216177#    ",
     "7471216177#    ",
     "7571216177#    ",
     "7671216177#    ",
     "7771216177#    ",
     "7871216177#    ",
     "7971216177#    ",
     "7A71216177#    ",
     "7B71216177#    ",
     "7C71216177#    ",
     "7D71216177#    ",
     "7*71216177#    ",
     "7601216177#    ",
     "7611216177#    ",
     "7621216177#    ",
     "7631216177#    ",
     "7641216177#    ",
     "7651216177#    ",
     "7661216177#    ",
     "7671216177#    ",
     "7681216177#    ",
     "7691216177#    ",
     "76A1216177#    ",
     "76B1216177#    ",
     "76C1216177#    ",
     "76D1216177#    ",
     "76*1216177#    ",
     "7670216177#    ",
     "7671216177#    ",
     "7672216177#    ",
     "7673216177#    ",
     "7674216177#    ",
     "7675216177#    ",
     "7676216177#    ",
     "7677216177#    ",
     "7678216177#    ",
     "7679216177#    ",
     "767A216177#    ",
     "767B216177#    ",
     "767C216177#    ",
     "767D216177#    ",
     "767*216177#    ",
     "7671016177#    ",
     "7671116177#    ",
     "7671216177#    ",
     "7671316177#    ",
     "7671416177#    ",
     "7671516177#    ",
     "7671616177#    ",
     "7671716177#    ",
     "7671816177#    ",
     "7671916177#    ",
     "7671A16177#    ",
     "7671B16177#    ",
     "7671C16177#    ",
     "7671D16177#    ",
     "7671*16177#    ",
     "7671206177#    ",
     "7671216177#    ",
     "7671226177#    ",
     "7671236177#    ",
     "7671246177#    ",
     "7671256177#    ",
     "7671266177#    ",
     "7671276177#    ",
     "7671286177#    ",
     "7671296177#    ",
     "76712A6177#    ",
     "76712B6177#    ",
     "76712C6177#    ",
     "76712D6177#    ",
     "76712*6177#    ",
     "7671210177#    ",
     "7671211177#    ",
     "7671212177#    ",
     "7671213177#    ",
     "7671214177#    ",
     "7671215177#    ",
     "7671216177#    ",
     "7671217177#    ",
     "7671218177#    ",
     "7671219177#    ",
     "767121A177#    ",
     "767121B177#    ",
     "767121C177#    ",
     "767121D177#    ",
     "767121*177#    ",
     "7671216077#    ",
     "7671216177#    ",
     "7671216277#    ",
     "7671216377#    ",
     "7671216477#    ",
     "7671216577#    ",
     "7671216677#    ",
     "7671216777#    ",
     "7671216877#    ",
     "7671216977#    ",
     "7671216A77#    ",
     "7671216B77#    ",
     "7671216C77#    ",
     "7671216D77#    ",
     "7671216*77#    ",
     "7671216107#    ",
     "7671216117#    ",
     "7671216127#    ",
     "7671216137#    ",
     "7671216147#    ",
     "7671216157#    ",
     "7671216167#    ",
     "7671216177#    ",
     "7671216187#    ",
     "7671216197#    ",
     "76712161A7#    ",
     "76712161B7#    ",
     "76712161C7#    ",
     "76712161D7#    ",
     "76712161*7#    ",
     "7671216170#    ",
     "7671216171#    ",
     "7671216172#    ",
     "7671216173#    ",
     "7671216174#    ",
     "7671216175#    ",
     "7671216176#    ",
     "7671216177#    ",
     "7671216178#    ",
     "7671216179#    ",
     "767121617A#    ",
     "767121617B#    ",
     "767121617C#    ",
     "767121617D#    ",
     "767121617*#    ",
     "00#            ",
     "01#            ",
     "02#            ",
     "03#            ",
     "04#            ",
     "05#            ",
     "06#            ",
     "07#            ",
     "08#            ",
     "09#            ",
     "0A#            ",
     "0B#            ",
     "0C#            ",
     "0D#            ",
     "0*#            ",
     "0#             ",
     "10#            ",
     "11#            ",
     "12#            ",
     "13#            ",
     "14#            ",
     "15#            ",
     "16#            ",
     "17#            ",
     "18#            ",
     "19#            ",
     "1A#            ",
     "1B#            ",
     "1C#            ",
     "1D#            ",
     "1*#            ",
     "1#             ",
     "20#            ",
     "21#            ",
     "22#            ",
     "23#            ",
     "24#            ",
     "25#            ",
     "26#            ",
     "27#            ",
     "28#            ",
     "29#            ",
     "2A#            ",
     "2B#            ",
     "2C#            ",
     "2D#            ",
     "2*#            ",
     "2#             ",
     "30#            ",
     "31#            ",
     "32#            ",
     "33#            ",
     "34#            ",
     "35#            ",
     "36#            ",
     "37#            ",
     "38#            ",
     "39#            ",
     "3A#            ",
     "3B#            ",
     "3C#            ",
     "3D#            ",
     "3*#            ",
     "3#             ",
     "40#            ",
     "41#            ",
     "42#            ",
     "43#            ",
     "44#            ",
     "45#            ",
     "46#            ",
     "47#            ",
     "48#            ",
     "49#            ",
     "4A#            ",
     "4B#            ",
     "4C#            ",
     "4D#            ",
     "4*#            ",
     "4#             ",
     "50#            ",
     "51#            ",
     "52#            ",
     "53#            ",
     "54#            ",
     "55#            ",
     "56#            ",
     "57#            ",
     "58#            ",
     "59#            ",
     "5A#            ",
     "5B#            ",
     "5C#            ",
     "5D#            ",
     "5*#            ",
     "5#             ",
     "60#            ",
     "61#            ",
     "62#            ",
     "63#            ",
     "64#            ",
     "65#            ",
     "66#            ",
     "67#            ",
     "68#            ",
     "69#            ",
     "6A#            ",
     "6B#            ",
     "6C#            ",
     "6D#            ",
     "6*#            ",
     "6#             ",
     "70#            ",
     "71#            ",
     "72#            ",
     "73#            ",
     "74#            ",
     "75#            ",
     "76#            ",
     "77#            ",
     "78#            ",
     "79#            ",
     "7A#            ",
     "7B#            ",
     "7C#            ",
     "7D#            ",
     "7*#            ",
     "7#             ",
     "80#            ",
     "81#            ",
     "82#            ",
     "83#            ",
     "84#            ",
     "85#            ",
     "86#            ",
     "87#            ",
     "88#            ",
     "89#            ",
     "8A#            ",
     "8B#            ",
     "8C#            ",
     "8D#            ",
     "8*#            ",
     "8#             ",
     "90#            ",
     "91#            ",
     "92#            ",
     "93#            ",
     "94#            ",
     "95#            ",
     "96#            ",
     "97#            ",
     "98#            ",
     "99#            ",
     "9A#            ",
     "9B#            ",
     "9C#            ",
     "9D#            ",
     "9*#            ",
     "9#             ",
     "A0#            ",
     "A1#            ",
     "A2#            ",
     "A3#            ",
     "A4#            ",
     "A5#            ",
     "A6#            ",
     "A7#            ",
     "A8#            ",
     "A9#            ",
     "AA#            ",
     "AB#            ",
     "AC#            ",
     "AD#            ",
     "A*#            ",
     "A#             ",
     "B0#            ",
     "B1#            ",
     "B2#            ",
     "B3#            ",
     "B4#            ",
     "B5#            ",
     "B6#            ",
     "B7#            ",
     "B8#            ",
     "B9#            ",
     "BA#            ",
     "BB#            ",
     "BC#            ",
     "BD#            ",
     "B*#            ",
     "B#             ",
     "C0#            ",
     "C1#            ",
     "C2#            ",
     "C3#            ",
     "C4#            ",
     "C5#            ",
     "C6#            ",
     "C7#            ",
     "C8#            ",
     "C9#            ",
     "CA#            ",
     "CB#            ",
     "CC#            ",
     "CD#            ",
     "C*#            ",
     "C#             ",
     "D0#            ",
     "D1#            ",
     "D2#            ",
     "D3#            ",
     "D4#            ",
     "D5#            ",
     "D6#            ",
     "D7#            ",
     "D8#            ",
     "D9#            ",
     "DA#            ",
     "DB#            ",
     "DC#            ",
     "DD#            ",
     "D*#            ",
     "D#             ",
     "*0#            ",
     "*1#            ",
     "*2#            ",
     "*3#            ",
     "*4#            ",
     "*5#            ",
     "*6#            ",
     "*7#            ",
     "*8#            ",
     "*9#            ",
     "*A#            ",
     "*B#            ",
     "*C#            ",
     "*D#            ",
     "**#            ",
     "*#             ",
     "7671216100#    ",
     "7671216101#    ",
     "7671216102#    ",
     "7671216103#    ",
     "7671216104#    ",
     "7671216105#    ",
     "7671216106#    ",
     "7671216107#    ",
     "7671216108#    ",
     "7671216109#    ",
     "767121610A#    ",
     "767121610B#    ",
     "767121610C#    ",
     "767121610D#    ",
     "767121610*#    ",
     "767121610#     ",
     "7671216110#    ",
     "7671216111#    ",
     "7671216112#    ",
     "7671216113#    ",
     "7671216114#    ",
     "7671216115#    ",
     "7671216116#    ",
     "7671216117#    ",
     "7671216118#    ",
     "7671216119#    ",
     "767121611A#    ",
     "767121611B#    ",
     "767121611C#    ",
     "767121611D#    ",
     "767121611*#    ",
     "767121611#     ",
     "7671216120#    ",
     "7671216121#    ",
     "7671216122#    ",
     "7671216123#    ",
     "7671216124#    ",
     "7671216125#    ",
     "7671216126#    ",
     "7671216127#    ",
     "7671216128#    ",
     "7671216129#    ",
     "767121612A#    ",
     "767121612B#    ",
     "767121612C#    ",
     "767121612D#    ",
     "767121612*#    ",
     "767121612#     ",
     "7671216130#    ",
     "7671216131#    ",
     "7671216132#    ",
     "7671216133#    ",
     "7671216134#    ",
     "7671216135#    ",
     "7671216136#    ",
     "7671216137#    ",
     "7671216138#    ",
     "7671216139#    ",
     "767121613A#    ",
     "767121613B#    ",
     "767121613C#    ",
     "767121613D#    ",
     "767121613*#    ",
     "767121613#     ",
     "7671216140#    ",
     "7671216141#    ",
     "7671216142#    ",
     "7671216143#    ",
     "7671216144#    ",
     "7671216145#    ",
     "7671216146#    ",
     "7671216147#    ",
     "7671216148#    ",
     "7671216149#    ",
     "767121614A#    ",
     "767121614B#    ",
     "767121614C#    ",
     "767121614D#    ",
     "767121614*#    ",
     "767121614#     ",
     "7671216150#    ",
     "7671216151#    ",
     "7671216152#    ",
     "7671216153#    ",
     "7671216154#    ",
     "7671216155#    ",
     "7671216156#    ",
     "7671216157#    ",
     "7671216158#    ",
     "7671216159#    ",
     "767121615A#    ",
     "767121615B#    ",
     "767121615C#    ",
     "767121615D#    ",
     "767121615*#    ",
     "767121615#     ",
     "7671216160#    ",
     "7671216161#    ",
     "7671216162#    ",
     "7671216163#    ",
     "7671216164#    ",
     "7671216165#    ",
     "7671216166#    ",
     "7671216167#    ",
     "7671216168#    ",
     "7671216169#    ",
     "767121616A#    ",
     "767121616B#    ",
     "767121616C#    ",
     "767121616D#    ",
     "767121616*#    ",
     "767121616#     ",
     "7671216170#    ",
     "7671216171#    ",
     "7671216172#    ",
     "7671216173#    ",
     "7671216174#    ",
     "7671216175#    ",
     "7671216176#    ",
     "7671216177#    ",
     "7671216178#    ",
     "7671216179#    ",
     "767121617A#    ",
     "767121617B#    ",
     "767121617C#    ",
     "767121617D#    ",
     "767121617*#    ",
     "767121617#     ",
     "7671216180#    ",
     "7671216181#    ",
     "7671216182#    ",
     "7671216183#    ",
     "7671216184#    ",
     "7671216185#    ",
     "7671216186#    ",
     "7671216187#    ",
     "7671216188#    ",
     "7671216189#    ",
     "767121618A#    ",
     "767121618B#    ",
     "767121618C#    ",
     "767121618D#    ",
     "767121618*#    ",
     "767121618#     ",
     "7671216190#    ",
     "7671216191#    ",
     "7671216192#    ",
     "7671216193#    ",
     "7671216194#    ",
     "7671216195#    ",
     "7671216196#    ",
     "7671216197#    ",
     "7671216198#    ",
     "7671216199#    ",
     "767121619A#    ",
     "767121619B#    ",
     "767121619C#    ",
     "767121619D#    ",
     "767121619*#    ",
     "767121619#     ",
     "76712161A0#    ",
     "76712161A1#    ",
     "76712161A2#    ",
     "76712161A3#    ",
     "76712161A4#    ",
     "76712161A5#    ",
     "76712161A6#    ",
     "76712161A7#    ",
     "76712161A8#    ",
     "76712161A9#    ",
     "76712161AA#    ",
     "76712161AB#    ",
     "76712161AC#    ",
     "76712161AD#    ",
     "76712161A*#    ",
     "76712161A#     ",
     "76712161B0#    ",
     "76712161B1#    ",
     "76712161B2#    ",
     "76712161B3#    ",
     "76712161B4#    ",
     "76712161B5#    ",
     "76712161B6#    ",
     "76712161B7#    ",
     "76712161B8#    ",
     "76712161B9#    ",
     "76712161BA#    ",
     "76712161BB#    ",
     "76712161BC#    ",
     "76712161BD#    ",
     "76712161B*#    ",
     "76712161B#     ",
     "76712161C0#    ",
     "76712161C1#    ",
     "76712161C2#    ",
     "76712161C3#    ",
     "76712161C4#    ",
     "76712161C5#    ",
     "76712161C6#    ",
     "76712161C7#    ",
     "76712161C8#    ",
     "76712161C9#    ",
     "76712161CA#    ",
     "76712161CB#    ",
     "76712161CC#    ",
     "76712161CD#    ",
     "76712161C*#    ",
     "76712161C#     ",
     "76712161D0#    ",
     "76712161D1#    ",
     "76712161D2#    ",
     "76712161D3#    ",
     "76712161D4#    ",
     "76712161D5#    ",
     "76712161D6#    ",
     "76712161D7#    ",
     "76712161D8#    ",
     "76712161D9#    ",
     "76712161DA#    ",
     "76712161DB#    ",
     "76712161DC#    ",
     "76712161DD#    ",
     "76712161D*#    ",
     "76712161D#     ",
     "76712161*0#    ",
     "76712161*1#    ",
     "76712161*2#    ",
     "76712161*3#    ",
     "76712161*4#    ",
     "76712161*5#    ",
     "76712161*6#    ",
     "76712161*7#    ",
     "76712161*8#    ",
     "76712161*9#    ",
     "76712161*A#    ",
     "76712161*B#    ",
     "76712161*C#    ",
     "76712161*D#    ",
     "76712161**#    ",
     "76712161*#     ",
     "07671216177#   ",
     "17671216177#   ",
     "27671216177#   ",
     "37671216177#   ",
     "47671216177#   ",
     "57671216177#   ",
     "67671216177#   ",
     "77671216177#   ",
     "87671216177#   ",
     "97671216177#   ",
     "A7671216177#   ",
     "B7671216177#   ",
     "C7671216177#   ",
     "D7671216177#   ",
     "*7671216177#   ",
     "70671216177#   ",
     "71671216177#   ",
     "72671216177#   ",
     "73671216177#   ",
     "74671216177#   ",
     "75671216177#   ",
     "76671216177#   ",
     "77671216177#   ",
     "78671216177#   ",
     "79671216177#   ",
     "7A671216177#   ",
     "7B671216177#   ",
     "7C671216177#   ",
     "7D671216177#   ",
     "7*671216177#   ",
     "76071216177#   ",
     "76171216177#   ",
     "76271216177#   ",
     "76371216177#   ",
     "76471216177#   ",
     "76571216177#   ",
     "76671216177#   ",
     "76771216177#   ",
     "76871216177#   ",
     "76971216177#   ",
     "76A71216177#   ",
     "76B71216177#   ",
     "76C71216177#   ",
     "76D71216177#   ",
     "76*71216177#   ",
     "76701216177#   ",
     "76711216177#   ",
     "76721216177#   ",
     "76731216177#   ",
     "76741216177#   ",
     "76751216177#   ",
     "76761216177#   ",
     "76771216177#   ",
     "76781216177#   ",
     "76791216177#   ",
     "767A1216177#   ",
     "767B1216177#   ",
     "767C1216177#   ",
     "767D1216177#   ",
     "767*1216177#   ",
     "76710216177#   ",
     "76711216177#   ",
     "76712216177#   ",
     "76713216177#   ",
     "76714216177#   ",
     "76715216177#   ",
     "76716216177#   ",
     "76717216177#   ",
     "76718216177#   ",
     "76719216177#   ",
     "7671A216177#   ",
     "7671B216177#   ",
     "7671C216177#   ",
     "7671D216177#   ",
     "7671*216177#   ",
     "76712016177#   ",
     "76712116177#   ",
     "76712216177#   ",
     "76712316177#   ",
     "76712416177#   ",
     "76712516177#   ",
     "76712616177#   ",
     "76712716177#   ",
     "76712816177#   ",
     "76712916177#   ",
     "76712A16177#   ",
     "76712B16177#   ",
     "76712C16177#   ",
     "76712D16177#   ",
     "76712*16177#   ",
     "76712106177#   ",
     "76712116177#   ",
     "76712126177#   ",
     "76712136177#   ",
     "76712146177#   ",
     "76712156177#   ",
     "76712166177#   ",
     "76712176177#   ",
     "76712186177#   ",
     "76712196177#   ",
     "767121A6177#   ",
     "767121B6177#   ",
     "767121C6177#   ",
     "767121D6177#   ",
     "767121*6177#   ",
     "76712160177#   ",
     "76712161177#   ",
     "76712162177#   ",
     "76712163177#   ",
     "76712164177#   ",
     "76712165177#   ",
     "76712166177#   ",
     "76712167177#   ",
     "76712168177#   ",
     "76712169177#   ",
     "7671216A177#   ",
     "7671216B177#   ",
     "7671216C177#   ",
     "7671216D177#   ",
     "7671216*177#   ",
     "76712161077#   ",
     "76712161177#   ",
     "76712161277#   ",
     "76712161377#   ",
     "76712161477#   ",
     "76712161577#   ",
     "76712161677#   ",
     "76712161777#   ",
     "76712161877#   ",
     "76712161977#   ",
     "76712161A77#   ",
     "76712161B77#   ",
     "76712161C77#   ",
     "76712161D77#   ",
     "76712161*77#   ",
     "76712161707#   ",
     "76712161717#   ",
     "76712161727#   ",
     "76712161737#   ",
     "76712161747#   ",
     "76712161757#   ",
     "76712161767#   ",
     "76712161777#   ",
     "76712161787#   ",
     "76712161797#   ",
     "767121617A7#   ",
     "767121617B7#   ",
     "767121617C7#   ",
     "767121617D7#   ",
     "767121617*7#   ",
     "76712161770#   ",
     "76712161771#   ",
     "76712161772#   ",
     "76712161773#   ",
     "76712161774#   ",
     "76712161775#   ",
     "76712161776#   ",
     "76712161777#   ",
     "76712161778#   ",
     "76712161779#   ",
     "7671216177A#   ",
     "7671216177B#   ",
     "7671216177C#   ",
     "7671216177D#   ",
     "7671216177*#   ",
     "671216177#     ",
     "771216177#     ",
     "761216177#     ",
     "767216177#     ",
     "767116177#     ",
     "767126177#     ",
     "767121177#     ",
     "767121677#     ",
     "767121617#     ",
     "767121617#     ",
     "#              ",
     "7#             ",
     "76#            ",
     "767#           ",
     "7671#          ",
     "76712#         ",
     "767121#        ",
     "7671216#       ",
     "76712161#      ",
     "767121617#     ",
     "7671216177#    ",
     "7671216177#    ",
     "671216177#     ",
     "71216177#      ",
     "1216177#       ",
     "216177#        ",
     "16177#         ",
     "6177#          ",
     "177#           ",
     "77#            ",
     "7#             ",
     "#              ",
     "767108088#     ",
     "767108088#     ",
     "767108088#     ",
     "767108088#     ",
     "767108088#     ",
     "767128088#     ",
     "767121088#     ",
     "767121688#     ",
     "767121618#     ",
     "767121617#     ",
     "7671216177#    ",
     "7671216177#    ",
     "7671216177#    ",
     "7671216177#    ",
     "7671216177#    ",
     "7671016177#    ",
     "7671086177#    ",
     "7671080177#    ",
     "7671080877#    ",
     "7671080887#    ",
     "767108088#     "
   ); 

end testbench_pkg;

package body testbench_pkg is
end testbench_pkg;
