library IEEE;
use IEEE.std_logic_1164.all;

package testbench_pkg is
   constant FILE_NAME : string := "chk_sim_sig_basic.txt";

   constant N_TEST_WORDS : integer := 48; 
   type t_test_words     is array (1 to N_TEST_WORDS) 
                                  of string(1 to 15);
   constant test_words : t_test_words :=
   ( 
     "767108088#     ",
     "1234567890*#   ",
     "767108088#     ",
     "234567890*#    ",
     "767108088#     ",
     "34567890*#     ",
     "767108088#     ",
     "4567890*#      ",
     "767108088#     ",
     "567890*#       ",
     "767108088#     ",
     "67890*#        ",
     "767108088#     ",
     "7890*#         ",
     "767108088#     ",
     "890*#          ",
     "767108088#     ",
     "90*#           ",
     "767108088#     ",
     "0*#            ",
     "767108088#     ",
     "*#             ",
     "767108088#     ",
     "#              ",
     "7671216177#    ",
     "1234567890*#   ",
     "7671216177#    ",
     "234567890*#    ",
     "7671216177#    ",
     "34567890*#     ",
     "7671216177#    ",
     "4567890*#      ",
     "7671216177#    ",
     "567890*#       ",
     "7671216177#    ",
     "67890*#        ",
     "7671216177#    ",
     "7890*#         ",
     "7671216177#    ",
     "890*#          ",
     "7671216177#    ",
     "90*#           ",
     "7671216177#    ",
     "0*#            ",
     "7671216177#    ",
     "*#             ",
     "7671216177#    ",
     "#              "
   ); 

end testbench_pkg;

package body testbench_pkg is
end testbench_pkg;
